
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY rom IS
    generic (n: integer:= 8); 
	PORT(

		clk : IN std_logic;
		we  : IN std_logic;
		address : IN  std_logic_vector(n-1 DOWNTO 0);
		datain  : IN  std_logic_vector(31 DOWNTO 0);
		dataout : OUT std_logic_vector(31 DOWNTO 0));
END ENTITY rom;

ARCHITECTURE syncroma OF rom IS
	--00000001000101101011001010000000
	--01000000010000011000000000001000
	TYPE rom_type IS ARRAY(0 TO 2**N -1) OF std_logic_vector(31 DOWNTO 0);
	SIGNAL rom : rom_type := (
        0=>"00000001000101101011001010000000",
	1=>"00000010001100100000000001000000",
	2=>"00000000001001000000000000000100",
	3=>"00000000000000000000000000000000",
	4=>"00000000000000000000000000000000",
	5=>"00000000000000000000000000000000",
	6=>"00000000000000000000000000000000",
	7=>"00000000000000000000000000000000",
	8=>"01000000010000011000000000001000",
	9=>"00000000000000000000000000000000",
	10=>"00000000000000000000000000000000",
	11=>"00000000000000000000000000000000",
	12=>"00000000000000000000000000000000",
	13=>"00000000000000000000000000000000",
	14=>"00000000000000000000000000000000",
	15=>"00000000000000000000000000000000",
	16=>"00101111010000001000000011000000",
	17=>"00000000000000000000000000000000",
	18=>"00000000000000000000000000000000",
	19=>"00000000000000000000000000000000",
	20=>"00000000000000000000000000000000",
	21=>"00000000000000000000000000000000",
	22=>"00000000000000000000000000000000",
	23=>"00000000000000000000000000000000",
	24=>"00011001010001101011001010000000",
	25=>"00101110001110000000000001010000",
	26=>"00000000000000000000000000000000",
	27=>"00000000000000000000000000000000",
	28=>"00000000000000000000000000000000",
	29=>"00000000000000000000000000000000",
	30=>"00000000000000000000000000000000",
	31=>"00000000000000000000000000000000",
	32=>"00100001010001100011010000000000",
	33=>"00101110001110001000000011010000",
	34=>"00000000000000000000000000000000",
	35=>"00000000000000000000000000000000",
	36=>"00000000000000000000000000000000",
	37=>"00000000000000000000000000000000",
	38=>"00000000000000000000000000000000",
	39=>"00000000000000000000000000000000",
	40=>"00101001000101101011001010000000",
	41=>"00101010010000000100000000000000", -- 51
	42=>"00101011001100100000000001000000", 
	43=>"00101100001001100000010000000000",
	44=>"00101110001100001000000011010000",
	45=>"00000000000000000000000000000000",
	46=>"00101111001000001000000011000000",
	47=>"01000000001000011000000000001000",
	48=>"00000000000000000000000000000000",
	49=>"00000000000000000000000000000000",
	50=>"00000000000000000000000000000000",
	51=>"00000000000000000000000000000000",
	52=>"00000000000000000000000000000000",
	53=>"00000000000000000000000000000000",
	54=>"00000000000000000000000000000000",
	55=>"00000000000000000000000000000000",
	56=>"00000000000000000000000000000000",
	57=>"00000000000000000000000000000000",
	58=>"00000000000000000000000000000000",
	59=>"00000000000000000000000000000000",
	60=>"00000000000000000000000000000000",
	61=>"00000000000000000000000000000000",
	62=>"00000000000000000000000000000000",
	63=>"00000000000000000000000000000000",
	64=>"10000000010100000100000000101000",
	65=>"00000000000000000000000000000000",
	66=>"00000000000000000000000000000000",
	67=>"00000000000000000000000000000000",
	68=>"00000000000000000000000000000000",
	69=>"00000000000000000000000000000000",
	70=>"00000000000000000000000000000000",
	71=>"00000000000000000000000000000000",
	72=>"01001001010101101011001010000000",
	73=>"01101110001110100000000001011000",
	74=>"00000000000000000000000000000000",
	75=>"00000000000000000000000000000000",
	76=>"00000000000000000000000000000000",
	77=>"00000000000000000000000000000000",
	78=>"00000000000000000000000000000000",
	79=>"00000000000000000000000000000000",
	80=>"01010001010101100011010000000000",
	81=>"01101110001110101000000011000000",
	82=>"00000000000000000000000000000000",
	83=>"00000000000000000000000000000000",
	84=>"00000000000000000000000000000000",
	85=>"00000000000000000000000000000000",
	86=>"00000000000000000000000000000000",
	87=>"00000000000000000000000000000000",
	88=>"01011001000101101011001010000000",
	89=>"01011010001100100000000000000000",
	90=>"01011011010100000100000001000000",
	91=>"01011100001001100000010000000000",
	92=>"01101110001100001000000011011000",
	93=>"00000000000000000000000000000000",
	94=>"00000000000000000000000000000000",
	95=>"00000000000000000000000000000000",
	96=>"01101111010100010000000011000000",
	97=>"00000000000000000000000000000000",
	98=>"00000000000000000000000000000000",
	99=>"00000000000000000000000000000000",
	100=>"00000000000000000000000000000000",
	101=>"00000000000000000000000000000000",
	102=>"00000000000000000000000000000000",
	103=>"00000000000000000000000000000000",
	104=>"00000000000000000000000000000000",
	105=>"00000000000000000000000000000000",
	106=>"00000000000000000000000000000000",
	107=>"00000000000000000000000000000000",
	108=>"00000000000000000000000000000000",
	109=>"00000000000000000000000000000000",
	110=>"01101111001000001000000011000000",
	111=>"10000000001000000100000000101000",
	112=>"00000000000000000000000000000000",
	113=>"00000000000000000000000000000000",
	114=>"00000000000000000000000000000000",
	115=>"00000000000000000000000000000000",
	116=>"00000000000000000000000000000000",
	117=>"00000000000000000000000000000000",
	118=>"00000000000000000000000000000000",
	119=>"00000000000000000000000000000000",
	120=>"00000000000000000000000000000000",
	121=>"00000000000000000000000000000000",
	122=>"00000000000000000000000000000000",
	123=>"00000000000000000000000000000000",
	124=>"00000000000000000000000000000000",
	125=>"00000000000000000000000000000000",
	126=>"00000000000000000000000000000000",
	127=>"00000000000000000000000000000000",
	128=>"00000000000000000000000000000000",
	129=>"10001010011101100000001000110000",
	130=>"10001010011101100000010000110000",
	131=>"10001010011101100000011000110000",
	132=>"10001010011101100000100000110000",
	133=>"10001010011101100000101000110000",
	134=>"10001010011101100000110000110000",
	135=>"10001010011101100000111000110000",
	136=>"10001010011101100001000000110000",
	137=>"10001010011101100000100000110000",
	138=>"11001100001100010000000101000000",
	139=>"11001100001110100000000000000000",
	140=>"00000000000000000000000000000000",
	141=>"00000000000000000000000000000000",
	142=>"00000000000000000000000000000000",
	143=>"00000000000000000000000000000000",
	144=>"00000000000000000000000000000000",
	145=>"00000000000000000000000000000000",
	146=>"00000000000000000000000000000000",
	147=>"00000000000000000000000000000000",
	148=>"00000000000000000000000000000000",
	149=>"00000000000000000000000000000000",
	150=>"00000000000000000000000000000000",
	151=>"00000000000000000000000000000000",
	152=>"00000000000000000000000000000000",
	153=>"00000000000000000000000000000000",
	154=>"00000000000000000000000000000000",
	155=>"00000000000000000000000000000000",
	156=>"00000000000000000000000000000000",
	157=>"00000000000000000000000000000000",
	158=>"00000000000000000000000000000000",
	159=>"00000000000000000000000000000000",
	160=>"10100001100000000100000000100000",
	161=>"10100010000101100000010000000000",
	162=>"10101001001100100000000000000000",
	163=>"00000000000000000000000000000000",
	164=>"00000000000000000000000000000000",
	165=>"00000000000000000000000000000000",
	166=>"00000000000000000000000000000000",
	167=>"00000000000000000000000000000000",
	168=>"00000000000000000000000000000000",
	169=>"00000000000000000000000000000001",
	170=>"00000000000000000000000000000000",
	171=>"00000000000000000000000000000000",
	172=>"00000000000000000000000000000000",
	173=>"00000000000000000000000000000000",
	174=>"00000000000000000000000000000000",
	175=>"00000000000000000000000000000000",
	176=>"00000000000000000000000000000000",
	177=>"00000000000000000000000000000000",
	178=>"00000000000000000000000000000000",
	179=>"00000000000000000000000000000000",
	180=>"00000000000000000000000000000000",
	181=>"00000000000000000000000000000000",
	182=>"00000000000000000000000000000000",
	183=>"00000000000000000000000000000000",
	184=>"00000000000000000000000000000000",
	185=>"00000000000000000000000000000000",
	186=>"00000000000000000000000000000000",
	187=>"00000000000000000000000000000000",
	188=>"00000000000000000000000000000000",
	189=>"00000000000000000000000000000000",
	190=>"00000000000000000000000000000000",
	191=>"00000000000000000000000000000000",
	192=>"11001010000001100010000000011000",
	193=>"11001010000001100010001000011000",
	194=>"11001010000001100010010000011000",
	195=>"11001010000001100010011000011000",
	196=>"11001010000001100010100000011000",
	197=>"11001010000001100010101000011000",
	198=>"11001010000001100010110000011000",
	199=>"11001010000001100010111000011000",
	200=>"11001010000001100011000000011000",
	201=>"00000000000000000000000000000000",
	202=>"11001100001100010000000101000000",
	203=>"11001100001110100000000000000000",
	204=>"00000000000000000000000000000001",
	205=>"00000000000000000000000000000000",
	206=>"00000000000000000000000000000000",
	207=>"00000000000000000000000000000000",
	208=>"00000000000000000000000000000000",
	209=>"00000000000000000000000000000000",
	210=>"00000000000000000000000000000000",
	211=>"00000000000000000000000000000000",
	212=>"00000000000000000000000000000000",
	213=>"00000000000000000000000000000000",
	214=>"00000000000000000000000000000000",
	215=>"00000000000000000000000000000000",
	216=>"00000000000000000000000000000000",
	217=>"00000000000000000000000000000000",
	218=>"00000000000000000000000000000000",
	219=>"00000000000000000000000000000000",
	220=>"00000000000000000000000000000000",
	221=>"00000000000000000000000000000000",
	222=>"00000000000000000000000000000000",
	223=>"00000000000000000000000000000000",
	224=>"00000000000000000000000000000000",
	225=>"00000000000000000000000000000000",
	226=>"00000000000000000000000000000000",
	227=>"00000000000000000000000000000000",
	228=>"00000000000000000000000000000000",
	229=>"00000000000000000000000000000000",
	230=>"00000000000000000000000000000000",
	231=>"00000000000000000000000000000000",
	232=>"00000000000000000000000000000000",
	233=>"00000000000000000000000000000000",
	234=>"00000000000000000000000000000000",
	235=>"00000000000000000000000000000000",
	236=>"00000000000000000000000000000000",
	237=>"00000000000000000000000000000000",
	238=>"00000000000000000000000000000000",
	239=>"00000000000000000000000000000000",
	240=>"00000000000000000000000000000000",
	241=>"00000000000000000000000000000000",
	242=>"00000000000000000000000000000000",
	243=>"00000000000000000000000000000000",
	244=>"00000000000000000000000000000000",
	245=>"00000000000000000000000000000000",
	246=>"00000000000000000000000000000000",
	247=>"00000000000000000000000000000000",
	248=>"00000000000000000000000000000000",
	249=>"00000000000000000000000000000000",
	250=>"00000000000000000000000000000000",
	251=>"00000000000000000000000000000000",
	252=>"00000000000000000000000000000000",
	253=>"00000000000000000000000000000000",
	254=>"00000000000000000000000000000000",
	255=>"00000000000000000000000000000010"
	        );
	
	BEGIN
		PROCESS(clk) IS
			BEGIN
				IF rising_edge(clk) THEN  
					IF we = '1' THEN
						rom(to_integer(unsigned(address))) <= datain;
					END IF;
				END IF;
		END PROCESS;
		dataout <= rom(to_integer(unsigned(address)));
END syncroma;